module Neuron(input clk, input rst);


endmodule
