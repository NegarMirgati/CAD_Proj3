module Controller(input clk, input rst, output acc_write, output ready);






endmodule
